module bullet_counter(); 

endmodule 