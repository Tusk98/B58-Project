// Possibly a file to keep track of where the bullet is onscreen and movement coordinates
module bullet_counter(); 

endmodule 