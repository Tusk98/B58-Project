module alien_counter();

endmodule