// Possibly a file to keep track of how many aliens there are on screen
module alien_counter();

endmodule